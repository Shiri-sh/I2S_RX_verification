interface i2s_if (input bit clk, input bit rstn);
    
    logic ws_i;
    logic sd_i;

endinterface