`include "uvm_macros.svh"


`include "cfg_pkg.sv"
`include "pcm_pkg.sv"
`include "i2s_pkg.sv"


`include "scoreboard.sv"
`include "env.sv" 
`include "virtual_sequence.sv"

`include "test_cfg_sterio.sv"
`include "test_cfg_mono_right.sv"
`include "test_cfg_mono_left.sv"
`include "test_enable.sv"

















