interface cfg_if ();
    logic clk;
    logic rstn;
    logic en;
    logic cfg_ch_single;
    logic cfg_ch_sel; 
endinterface